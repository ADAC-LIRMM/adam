/*
 * Copyright 2025 LIRMM
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

interface ADAM_STREAM #(
    parameter type T = logic
);

    T     data;
    logic valid;
    logic ready;

    modport Master (
        output data,
        output valid,
        input  ready
    );

    modport Slave (
        input  data,
        input  valid,
        output ready
    );

endinterface

interface ADAM_STREAM_DV #(
    parameter type T = logic
) (
    input logic clk
);

    T     data;
    logic valid;
    logic ready;
    
    modport Master (
        output data,
        output valid,
        input  ready
    );

    modport Slave (
        input  data,
        input  valid,
        output ready
    );

endinterface