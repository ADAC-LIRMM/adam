/*
 * Copyright 2025 LIRMM
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

module adam_clk_gate (
    ADAM_SEQ.Slave  slv,
    ADAM_SEQ.Master mst,

    input  logic enable
);

    logic ctrl;

    always_latch begin
        if (slv.clk == 0) ctrl <= enable | slv.rst;
    end

    assign mst.rst = slv.rst;
    assign mst.clk = slv.clk & ctrl;

endmodule
