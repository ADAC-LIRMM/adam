/*
 * Copyright 2025 LIRMM
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

`timescale 1ns/1ps
`include "adam/macros_bhv.svh"

module adam_seq_bhv #(
    `ADAM_BHV_CFG_PARAMS
) (
    ADAM_SEQ.Master seq
);

    initial begin
        seq.clk <= 1;
        forever #(CLK_PERIOD/2) seq.clk <= ~seq.clk;
    end

    initial begin
        seq.rst <= 1;
        repeat (RST_CYCLES) @(posedge seq.clk);
        seq.rst <= #TA 0;
    end

endmodule