`timescale 1ns/1ps
`include "adam/macros_bhv.svh"
`include "vunit_defines.svh"

module adam_tb;
    import adam_jtag_mst_bhv::*;

    `ADAM_BHV_CFG_LOCALPARAMS;
    
    localparam integer LPMEM_SIZE = 1024;

    localparam integer MEM_SIZE [NO_MEMS+1] = 
        '{32768, 32768, 32768, 0};

    // seq and pause ==========================================================

    ADAM_SEQ lsdom_seq ();
    ADAM_SEQ hsdom_seq ();

    ADAM_PAUSE lsdom_pause_ext ();

    adam_seq_bhv #(
        `ADAM_BHV_CFG_PARAMS_MAP
    ) lsdom_adam_seq_bhv (
        .seq (lsdom_seq)
    );

    adam_seq_bhv #(
        `ADAM_BHV_CFG_PARAMS_MAP
    ) hsdom_adam_seq_bhv (
        .seq (hsdom_seq)
    );

    `ADAM_PAUSE_MST_TIE_ON(lsdom_pause_ext);

    // lpmem ==================================================================

    logic        lsdom_lpmem_rst;
    ADAM_SEQ     lsdom_lpmem_seq ();
    ADAM_PAUSE   lsdom_lpmem_pause ();
    `ADAM_AXIL_I lsdom_lpmem_axil ();

    logic  lsdom_lpmem_req;
    ADDR_T lsdom_lpmem_addr;
    logic  lsdom_lpmem_we;
    STRB_T lsdom_lpmem_be;
    DATA_T lsdom_lpmem_wdata;
    DATA_T lsdom_lpmem_rdata;

    assign lsdom_lpmem_seq.clk = lsdom_seq.clk;
    assign lsdom_lpmem_seq.rst = lsdom_seq.rst || lsdom_lpmem_rst;

    if (EN_LPMEM) begin
        adam_axil_to_mem #(
            `ADAM_CFG_PARAMS_MAP
        ) adam_axil_to_mem (
            .seq   (lsdom_lpmem_seq),
            .pause (lsdom_lpmem_pause),

            .axil (lsdom_lpmem_axil),

            .mem_req   (lsdom_lpmem_req),
            .mem_addr  (lsdom_lpmem_addr),
            .mem_we    (lsdom_lpmem_we),
            .mem_be    (lsdom_lpmem_be),
            .mem_wdata (lsdom_lpmem_wdata),
            .mem_rdata (lsdom_lpmem_rdata)
        );

        adam_mem #(
            `ADAM_CFG_PARAMS_MAP,

            .SIZE (LPMEM_SIZE)
        ) adam_mem (
            .seq (lsdom_lpmem_seq),

            .req   (lsdom_lpmem_req),
            .addr  (lsdom_lpmem_addr),
            .we    (lsdom_lpmem_we),
            .be    (lsdom_lpmem_be),
            .wdata (lsdom_lpmem_wdata),
            .rdata (lsdom_lpmem_rdata)
        );
    end
    else begin
        // TODO: tie off
    end

    // mem ====================================================================
    
    logic        hsdom_mem_rst   [NO_MEMS+1];
    ADAM_SEQ     hsdom_mem_seq   [NO_MEMS+1] ();
    ADAM_PAUSE   hsdom_mem_pause [NO_MEMS+1] ();
    `ADAM_AXIL_I hsdom_mem_axil  [NO_MEMS+1] ();
    
    logic  hsdom_mem_req   [NO_MEMS+1];
    ADDR_T hsdom_mem_addr  [NO_MEMS+1];
    logic  hsdom_mem_we    [NO_MEMS+1];
    STRB_T hsdom_mem_be    [NO_MEMS+1];
    DATA_T hsdom_mem_wdata [NO_MEMS+1];
    DATA_T hsdom_mem_rdata [NO_MEMS+1];

    for (genvar i = 0; i < NO_MEMS; i++) begin
        assign hsdom_mem_seq[i].clk = lsdom_seq.clk;
        assign hsdom_mem_seq[i].rst = lsdom_seq.rst || hsdom_mem_rst[i];

        adam_axil_to_mem #(
            `ADAM_CFG_PARAMS_MAP
        ) adam_axil_to_mem (
            .seq   (hsdom_mem_seq[i]),
            .pause (hsdom_mem_pause[i]),

            .axil (hsdom_mem_axil[i]),

            .mem_req   (hsdom_mem_req[i]),
            .mem_addr  (hsdom_mem_addr[i]),
            .mem_we    (hsdom_mem_we[i]),
            .mem_be    (hsdom_mem_be[i]),
            .mem_wdata (hsdom_mem_wdata[i]),
            .mem_rdata (hsdom_mem_rdata[i])
        );
    end

    // sensemark #(
    //     `ADAM_CFG_PARAMS_MAP
    // ) sensemark (
    //     .seq (hsdom_mem_seq[0]),

    //     .req   (hsdom_mem_req[0]),
    //     .addr  (hsdom_mem_addr[0]),
    //     .we    (hsdom_mem_we[0]),
    //     .be    (hsdom_mem_be[0]),
    //     .wdata (hsdom_mem_wdata[0]),
    //     .rdata (hsdom_mem_rdata[0])
    // );

    for (genvar i = 0; i < NO_MEMS; i++) begin
        adam_mem #(
            `ADAM_CFG_PARAMS_MAP,

            .SIZE (MEM_SIZE[i])
        ) adam_mem (
            .seq (hsdom_mem_seq[i]),

            .req   (hsdom_mem_req[i]),
            .addr  (hsdom_mem_addr[i]),
            .we    (hsdom_mem_we[i]),
            .be    (hsdom_mem_be[i]),
            .wdata (hsdom_mem_wdata[i]),
            .rdata (hsdom_mem_rdata[i])
        );
    end
    
    // lspa io ================================================================

    ADAM_IO     lspa_gpio_io   [NO_LSPA_GPIOS*GPIO_WIDTH+1] ();
    logic [1:0] lspa_gpio_func [NO_LSPA_GPIOS*GPIO_WIDTH+1];

    ADAM_IO lspa_spi_sclk [NO_LSPA_SPIS+1] ();
    ADAM_IO lspa_spi_mosi [NO_LSPA_SPIS+1] ();
    ADAM_IO lspa_spi_miso [NO_LSPA_SPIS+1] ();
    ADAM_IO lspa_spi_ss_n [NO_LSPA_SPIS+1] ();

    ADAM_IO lspa_uart_tx [NO_LSPA_UARTS+1] ();
    ADAM_IO lspa_uart_rx [NO_LSPA_UARTS+1] ();

    for (genvar i = 0; i < NO_LSPA_GPIOS; i++) begin
        `ADAM_IO_SLV_TIE_OFF(lspa_gpio_io[i]);
    end
    for (genvar i = 0; i < NO_LSPA_SPIS; i++) begin
        `ADAM_IO_SLV_TIE_OFF(lspa_spi_sclk[i]);
        `ADAM_IO_SLV_TIE_OFF(lspa_spi_mosi[i]);
        `ADAM_IO_SLV_TIE_OFF(lspa_spi_miso[i]);
        `ADAM_IO_SLV_TIE_OFF(lspa_spi_ss_n[i]);
    end
    for (genvar i = 0; i < NO_LSPA_UARTS; i++) begin
        `ADAM_IO_SLV_TIE_OFF(lspa_uart_tx[i]);
        `ADAM_IO_SLV_TIE_OFF(lspa_uart_rx[i]);
    end

    // lspb io ================================================================

    ADAM_IO     lspb_gpio_io   [NO_LSPB_GPIOS*GPIO_WIDTH+1] ();
    logic [1:0] lspb_gpio_func [NO_LSPB_GPIOS*GPIO_WIDTH+1];

    ADAM_IO lspb_spi_sclk [NO_LSPB_SPIS+1] ();
    ADAM_IO lspb_spi_mosi [NO_LSPB_SPIS+1] ();
    ADAM_IO lspb_spi_miso [NO_LSPB_SPIS+1] ();
    ADAM_IO lspb_spi_ss_n [NO_LSPB_SPIS+1] ();

    ADAM_IO lspb_uart_tx [NO_LSPB_UARTS+1] ();
    ADAM_IO lspb_uart_rx [NO_LSPB_UARTS+1] ();

    for (genvar i = 0; i < NO_LSPB_GPIOS; i++) begin
        `ADAM_IO_SLV_TIE_OFF(lspb_gpio_io[i]);
    end
    for (genvar i = 0; i < NO_LSPB_SPIS; i++) begin
        `ADAM_IO_SLV_TIE_OFF(lspb_spi_sclk[i]);
        `ADAM_IO_SLV_TIE_OFF(lspb_spi_mosi[i]);
        `ADAM_IO_SLV_TIE_OFF(lspb_spi_miso[i]);
        `ADAM_IO_SLV_TIE_OFF(lspb_spi_ss_n[i]);
    end
    for (genvar i = 0; i < NO_LSPB_UARTS; i++) begin
        `ADAM_IO_SLV_TIE_OFF(lspb_uart_tx[i]);
        `ADAM_IO_SLV_TIE_OFF(lspb_uart_rx[i]);
    end

    // debug ==================================================================

    ADAM_JTAG jtag ();

    adam_jtag_mst_bhv #(
        `ADAM_BHV_CFG_PARAMS_MAP
    ) jtag_bhv;

    // dut ====================================================================

    adam #(
        `ADAM_CFG_PARAMS_MAP
    ) dut (
        .lsdom_seq (lsdom_seq),

        .lsdom_pause_ext  (lsdom_pause_ext),

        .lsdom_lpmem_rst   (lsdom_lpmem_rst),
        .lsdom_lpmem_pause (lsdom_lpmem_pause),
        .lsdom_lpmem_axil  (lsdom_lpmem_axil),

        .hsdom_seq       (hsdom_seq),

        .hsdom_mem_rst   (hsdom_mem_rst),
        .hsdom_mem_pause (hsdom_mem_pause),
        .hsdom_mem_axil  (hsdom_mem_axil),
        
        .jtag (jtag),

        .lspa_gpio_io   (lspa_gpio_io),
        .lspa_gpio_func (lspa_gpio_func),

        .lspa_spi_sclk (lspa_spi_sclk),
        .lspa_spi_mosi (lspa_spi_mosi),
        .lspa_spi_miso (lspa_spi_miso),
        .lspa_spi_ss_n (lspa_spi_ss_n),

        .lspa_uart_tx (lspa_uart_tx),
        .lspa_uart_rx (lspa_uart_rx),
        
        .lspb_gpio_io   (lspb_gpio_io),
        .lspb_gpio_func (lspb_gpio_func),

        .lspb_spi_sclk (lspb_spi_sclk),
        .lspb_spi_mosi (lspb_spi_mosi),
        .lspb_spi_miso (lspb_spi_miso),
        .lspb_spi_ss_n (lspb_spi_ss_n),

        .lspb_uart_tx (lspb_uart_tx),
        .lspb_uart_rx (lspb_uart_rx)
    );

    // test ===================================================================

    localparam W_IR = 5;
    
    localparam IDLE  = 1;
    localparam ABITS = 7;
    
    localparam A_IDCODE = 'h01;
    localparam A_DTMCS  = 'h10;
    localparam A_DMI    = 'h11;

    localparam W_IDCODE = 32;
    localparam W_DTMCS  = 32;
    localparam W_DMI    = ABITS+34;

    localparam A_DMCONTROL  = 'h10;
    localparam A_DMSTATUS   = 'h11;
    localparam A_SBCS       = 'h38;
    localparam A_SBADDRESS0 = 'h39;
    localparam A_SBDATA0    = 'h3C;

    typedef logic[ABITS-1:0] dmaddr_t;
    typedef logic[31:0]      dmdata_t;

    `TEST_SUITE begin
        `TEST_CASE("minimal") begin
            jtag_bhv = new(jtag);
            #10us;
        end

        `TEST_CASE("debug") begin
            ADDR_T  addr;
            DATA_T  wdata;
            DATA_T  rdata;

            addr  = 32'h0100_0000;
            wdata = 32'hDEAD_BEEF;

            jtag_bhv = new(jtag);

            if (EN_DEBUG) begin
                dtm_init();
                dm_init();          
                dm_select('d1); // HART 1 aka CPU0
                dm_halt();
                
                if (EN_BOOTSTRAP_MEM0) begin
                    dm_sb_write(addr, wdata);
                    dm_sb_read(addr, rdata);
                    assert (rdata == wdata);
                end

                dm_resume();
            end
        end
    end

    initial begin
        #1000us $error("timeout");
    end

    task dtm_init();
        logic [W_IDCODE-1:0] idcode;
        logic [W_DTMCS-1:0] dtmcs;

        $display("dtm_init start");

        jtag_bhv.reset();
        jtag_bhv.tap_reset();

        jtag_bhv.tap_reg_read(A_IDCODE, W_IR, idcode, W_IDCODE);
        assert(idcode == DEBUG_IDCODE);

        jtag_bhv.tap_reg_read(A_DTMCS, W_IR, dtmcs, W_DTMCS);
        assert(dtmcs[9:4] == ABITS);
        assert(dtmcs[14:12] == IDLE);

        $display("dtm_init end");
    endtask

    task dm_init();
        $display("dm_init start");
        
        dm_write(A_DMCONTROL, '1); // set dmactive

        $display("dm_init end");
    endtask

    task dm_select(
        input [19:0] hartsel
    );
        dmdata_t dmcontrol;

        $display("dm_select start");

        dm_read(A_DMCONTROL, dmcontrol);

        dmcontrol[25:6] = {hartsel[ 9: 0], hartsel[19:10]};
        dm_write(A_DMCONTROL, dmcontrol);

        dm_read(A_DMCONTROL, dmcontrol);
        assert(dmcontrol[25:6] == {hartsel[ 9: 0], hartsel[19:10]});

        $display("dm_select end");
    endtask

    task dm_halt();
        dmdata_t dmcontrol;
        dmdata_t dmstatus;

        $display("dm_halt start");

        dm_read(A_DMCONTROL, dmcontrol);

        // set haltreq
        dmcontrol[31] = '1;
        dm_write(A_DMCONTROL, dmcontrol);

        // wait of allhalted
        do begin
            dm_read(A_DMSTATUS, dmstatus);
        end while (!dmstatus[9]);

        // clear haltreq
        dmcontrol[31] = '0;
        dm_write(A_DMCONTROL, dmcontrol);

        $display("dm_halt end");
    endtask

    task dm_resume();
        dmdata_t dmcontrol;
        dmdata_t dmstatus;

        $display("dm_resume start");

        // set resumereq
        dm_read(A_DMCONTROL, dmcontrol);
        dmcontrol[30] = '1;
        dm_write(A_DMCONTROL, dmcontrol);

        // wait allresumeack
        do begin
            dm_read(A_DMSTATUS, dmstatus);
        end while (!dmstatus[17]);

        // clear resumereq
        dmcontrol[30] = '0;
        dm_write(A_DMCONTROL, dmcontrol);  

        $display("dm_resume end");      
    endtask

    task dm_sb_write(
        input ADDR_T addr,
        input DATA_T data
    );
        dmdata_t sbcs;

        dm_bus_wait();

        // clear sbreadonaddr
        dm_read(A_SBCS, sbcs);
        sbcs[20] = '0;
        dm_write(A_SBCS, sbcs);

        // write to address0
        dm_write(A_SBADDRESS0, addr);

        // write to sbdata0
        dm_write(A_SBDATA0, data);

        dm_bus_wait();
    endtask

    task dm_sb_read(
        input  ADDR_T addr,
        output DATA_T data
    );
        dmdata_t sbcs;

        dm_bus_wait();

        // set sbreadonaddr
        dm_read(A_SBCS, sbcs);
        sbcs[20] = '1; 
        dm_write(A_SBCS, sbcs);

        // write to address0
        dm_write(A_SBADDRESS0, addr);

        dm_bus_wait();

        // write to sbdata0
        dm_read(A_SBDATA0, data);
    endtask

    task dm_bus_wait();
        dmdata_t sbcs;

        // wait sbbusy
        do begin
            dm_read(A_SBCS, sbcs);
        end while (sbcs[21]);
    endtask

    task dm_read(
        input  dmaddr_t addr,
        output dmdata_t data 
    );
        logic [W_DMI-1:0] dmi;
        
        dmi[ABITS+33:34] = addr;
        dmi[33:2] = '0; 
        dmi[1:0] = 'd1;
        jtag_bhv.tap_reg_write(A_DMI, W_IR, dmi, W_DMI);
        
        repeat (IDLE-1) jtag_bhv.tap_nop();
        
        jtag_bhv.tap_reg_read(A_DMI, W_IR, dmi, W_DMI);
        assert(dmi[1:0] == '0);
        data = dmi[33:2];
    endtask

    task dm_write(
        input dmaddr_t addr,
        input dmdata_t data 
    );
        logic [31:0] idcode;
        logic [ABITS+33:0] dmi;
        
        dmi[ABITS+33:34] = addr;
        dmi[33:2] = data; 
        dmi[1:0] = 'd2;
        jtag_bhv.tap_reg_write(A_DMI, W_IR, dmi, W_DMI);
        
        repeat (IDLE-1) jtag_bhv.tap_nop();
        
        jtag_bhv.tap_reg_read (A_DMI, W_IR, dmi, W_DMI);
        assert(dmi[1:0] == 0); // check if op is 0
    endtask

endmodule
