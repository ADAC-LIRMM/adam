/*
 * Copyright 2025 LIRMM
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

interface ADAM_JTAG;

    logic trst_n;
    logic tck;
    logic tms;
    logic tdi;
    logic tdo;

    modport Master (
        output trst_n,
        output tck,
        output tms,
        output tdi,
        input  tdo
    );

    modport Slave (
        input  trst_n,
        input  tck,
        input  tms,
        input  tdi,
        output tdo
    );

endinterface